library verilog;
use verilog.vl_types.all;
entity full_test is
end full_test;
